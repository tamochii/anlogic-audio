`timescale 1ns/1ns

module es8388_config(
    input        clk     ,                  // ʱ���ź�
    input        rst_n   ,                  // ��λ�ź�
    
	 input  [1:0] volume ,                  //������������
	 
    output       aud_scl ,                  // es8388��SCLʱ��
    inout        aud_sda                    // es8388��SDA�ź�
);

//parameter define
parameter   SLAVE_ADDR = 7'h10         ;    // es8388������ַ
parameter   WL         = 6'd32         ;    // word length��Ƶ�ֳ���������
parameter   BIT_CTRL   = 1'b0          ;    // �ֵ�ַλ���Ʋ���(16b/8b)
parameter   CLK_FREQ   = 26'd50_000_000;    // i2c_driģ�������ʱ��Ƶ��(CLK_FREQ)
parameter   I2C_FREQ   = 18'd250_000   ;    // I2C��SCLʱ��Ƶ��

//wire define
wire        clk_i2c   ;                     // i2c�Ĳ���ʱ��
wire        i2c_exec  ;                     // i2c��������
wire        i2c_done  ;                     // i2c����������־
wire        cfg_done  ;                     // es8388������ɱ�־
wire [15:0] reg_data  ;                     // es8388��Ҫ���õļĴ�������ַ�����ݣ�

//*****************************************************
//**                    main code
//*****************************************************

//����es8388�ļĴ���
i2c_reg_cfg #(
    .WL             (WL       )             // word length��Ƶ�ֳ���������
) u_i2c_reg_cfg(  
    .clk            (clk_i2c  ),            // i2c_reg_cfg����ʱ��
    .rst_n          (rst_n    ),            // ��λ�ź�
  
    .i2c_exec       (i2c_exec ),            // I2C����ִ���ź�
    .i2c_data       (reg_data ),            // �Ĵ������ݣ�7λ��ַ+9λ���ݣ�
    
	 .volume         (volume),              //������������
	 
    .i2c_done       (i2c_done ),            // I2Cһ�β�����ɵı�־�ź�            
    .cfg_done       (cfg_done )             // es8388�������
);

//����IICЭ��
i2c_dri #(
    .SLAVE_ADDR     (SLAVE_ADDR),           // slave address�ӻ���ַ���Ŵ˴������������
    .CLK_FREQ       (CLK_FREQ  ),           // i2c_driģ�������ʱ��Ƶ��(CLK_FREQ)
    .I2C_FREQ       (I2C_FREQ  )            // I2C��SCLʱ��Ƶ��
) u_i2c_dri(  
    .clk            (clk       ),           // i2c_driģ�������ʱ��(CLK_FREQ)
    .rst_n          (rst_n     ),           // ��λ�ź�
  
    .i2c_exec       (i2c_exec  ),           // I2C����ִ���ź�
    .bit_ctrl       (BIT_CTRL  ),           // ������ַλ����(16b/8b)
    .i2c_rh_wl      (1'b0      ),           // I2C��д�����ź�
    .i2c_addr       (reg_data[15:8]),       // I2C�����ֵ�ַ
    .i2c_data_w     (reg_data[ 7:0]),       // I2CҪд������
      
    .i2c_data_r     (),                     // I2C����������
    .i2c_done       (i2c_done  ),           // I2Cһ�β������
      
    .scl            (aud_scl   ),           // I2C��SCLʱ���ź�
    .sda            (aud_sda   ),           // I2C��SDA�ź�
    .dri_clk        (clk_i2c   )            // I2C����ʱ��
);

endmodule 